module test1(
	input a,
	input b,
	output result
	);
	
	assign result = a|b;
	
endmodule